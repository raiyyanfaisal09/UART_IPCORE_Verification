`define ADDR 3
`define DATA 8
