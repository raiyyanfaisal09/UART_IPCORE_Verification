class wr_seqs extends uvm_sequence #(write_xtn);
`uvm_object_utils(wr_seqs)




endclass
